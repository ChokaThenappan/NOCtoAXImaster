function [1:0] get_msg_type;
    ;
    
endfunction